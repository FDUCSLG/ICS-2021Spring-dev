`include "defs.sv"
